entity tb is
  generic (
    genInt : integer := 42;
    genStr : string := "default string"
  );
end entity;
