
entity ent is
end entity ent;

architecture behavioral of ent is
begin
end architecture behavioral;

