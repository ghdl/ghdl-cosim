library ieee;
context ieee.ieee_std_context;

package vffi_user is

  function reverseBitsInBytes (datain : std_logic_vector(0 to 127)) return std_logic_vector;

end vffi_user;
